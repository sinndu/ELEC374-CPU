// Testbench for SHL instruction
`timescale 1ns/10ps
module DataPath_tb_rol;
    reg [3:0] reg_select;
    reg PCout, Zlowout, MDRout, Rout;
    reg MARin, Zin, PCin, MDRin, IRin, Yin;
    reg Read, Rin;
    reg Clock, clear;
    reg [31:0] Mdatain;
    parameter   Default = 4'b0000, Reg_load1a = 4'b0001, Reg_load1b = 4'b0010, Reg_load2a = 4'b0011,
                Reg_load2b = 4'b0100, Reg_load3a = 4'b0101, Reg_load3b = 4'b0110, T0 = 4'b0111,
                T1 = 4'b1000, T2 = 4'b1001, T3 = 4'b1010, T4 = 4'b1011, T5 = 4'b1100, done = 4'b1101;
    reg [3:0] Present_state = Default;

    parameter   ADD = 4'b0000, SUB = 4'b0001, AND = 4'b0010, OR = 4'b011, NEG = 4'b0100, NOT = 4'b0101, 
                SHR = 4'b0110, SHRA = 4'b0111, SHL = 4'b1000, ROR = 4'b1001, ROL = 4'b1010,
                MUL = 4'b1011, DIV = 4'b1100, IncPC = 4'b1101, NONE = 4'b1110;
    reg [3:0] ALU_operation = NONE;

datapath DUT(

    .clock(Clock), .clear(clear),
    .in_memory_data(Mdatain),
    .PCin(PCin), .PCout(PCout), 		
    .IRin(IRin),
    .ZLowout(Zlowout), 
    .MARin(MARin), .MDRin(MDRin), .MDRout(MDRout), .read(Read),
    .Rin(Rin), .Rout(Rout), 
    .Yin(Yin), .Zin(Zin),
    .ALU_operation(ALU_operation), 
    .reg_select(reg_select)

);

// add test logic here
initial
    begin
		Clock = 0;
		forever #10 Clock = ~ Clock;
end

initial 
	begin
		clear = 1;
		#25;
		clear = 0;
end

always @(posedge Clock) // finite state machine; if clock rising-edge
    begin
        case (Present_state)
            Default : Present_state = Reg_load1a;
            Reg_load1a : Present_state = Reg_load1b;
            Reg_load1b : Present_state = Reg_load2a;
            Reg_load2a : Present_state = Reg_load2b;
            Reg_load2b : Present_state = Reg_load3a;
            Reg_load3a : Present_state = Reg_load3b;
            Reg_load3b : Present_state = T0;
            T0 : Present_state = T1;
            T1 : Present_state = T2;
            T2 : Present_state = T3;
            T3 : Present_state = T4;
            T4 : Present_state = T5;
				T5 : Present_state = done;
        endcase
    end

always @(negedge Clock) // do the required job in each state
    begin
    //clear all signals before switch case
    PCout <= 0; Zlowout <= 0; MDRout <= 0; Rout <= 0;
    MARin <= 0; Zin <= 0; PCin <= 0; MDRin <= 0;
    IRin <= 0; Yin <= 0; Read <= 0;
    Rin <= 0; ALU_operation <= NONE;

        case (Present_state) // assert the required signals in each clock cycle
            Default: begin
                        PCout = 0; Zlowout = 0; MDRout = 0; // initialize the signals
                        Rout = 0; MARin = 0; Zin = 0;
                        PCin = 0; MDRin = 0; IRin = 0; Yin = 0;
                        Read = 0; ALU_operation = NONE;
                        Rin = 0; Mdatain = 32'h00000000;
            end
            Reg_load1a: begin
								
                        Mdatain <= 32'hFFFFFFFE;
                        Read <= 1; MDRin <= 1; 
            end
            Reg_load1b: begin
                        MDRout <= 1; reg_select <= 0; Rin <= 1;
                        // initialize R0 with the value 0xFFFF
            end
            Reg_load2a: begin
                        Mdatain <= 32'h00000001;
                        Read <= 1; MDRin <= 1;
            end
            Reg_load2b: begin
                        MDRout <= 1; reg_select <= 4; Rin <= 1;
                        // initialize R4 with the value 0x1
            end
            Reg_load3a: begin
                        Mdatain <= 32'h00000067;
                        Read <= 1; MDRin <= 1;
                        
            end
            Reg_load3b: begin
                        MDRout <= 1; reg_select <= 2; Rin <= 1;
                        // initialize R7 with the value 0x67
            end
            T0: begin // see if you need to de-assert these signals
                        PCout <= 1; MARin <= 1; ALU_operation <= IncPC; Zin <= 1;
            end
            T1: begin
                        Zlowout <= 1; PCin <= 1; Read <= 1; MDRin <= 1;
                        Mdatain <= 32'h112B0000; // opcode
            end
            T2: begin
                        MDRout <= 1; IRin <= 1;
            end
            T3: begin
                        reg_select <= 0; Rout <= 1; Yin <= 1;
            end
            T4: begin
                        reg_select <= 4; Rout <= 1; ALU_operation <= ROL; Zin <= 1;
            end
            T5: begin
                        Zlowout <= 1; reg_select <= 7; Rin <= 1;
            end
        endcase
    end
	 
always @(negedge Clock) begin 
	case (Present_state)
		T0: begin
			$display(
				"T0 @ %0t | PC=%0d MAR=%h MDR=%h IR=%h ALU_op=%0d Zlow=%0d reg_select=%b  R7=%h R0=%h R4=%h Y=%h Bus=%h",
				$time, DUT.PC.storage, DUT.MAR.storage, DUT.MDR.MDR_Reg.storage, DUT.IR.storage, ALU_operation, DUT.RZlow.storage, DUT.reg_decode, DUT.R7.storage, DUT.R5.storage, DUT.R6.storage, DUT.RY.storage, DUT.bus.q,
			);
		end
		T1: begin
			$display(
				"T1 @ %0t | PC=%0d MAR=%h MDR=%h IR=%h ALU_op=%0d Zlow=%0d reg_select=%b  R7=%h R0=%h R4=%h Y=%h Bus=%h",
				$time, DUT.PC.storage, DUT.MAR.storage, DUT.MDR.MDR_Reg.storage, DUT.IR.storage, ALU_operation, DUT.RZlow.storage, DUT.reg_decode, DUT.R7.storage, DUT.R0.storage, DUT.R4.storage, DUT.RY.storage, DUT.bus.q,
			);
		end
		T2: begin
			$display(
				"T2 @ %0t | PC=%0d MAR=%h MDR=%h IR=%h ALU_op=%0d Zlow=%0d reg_select=%b  R7=%h R0=%h R4=%h Y=%h Bus=%h",
				$time, DUT.PC.storage, DUT.MAR.storage, DUT.MDR.MDR_Reg.storage, DUT.IR.storage, ALU_operation, DUT.RZlow.storage, DUT.reg_decode, DUT.R7.storage, DUT.R0.storage, DUT.R4.storage, DUT.RY.storage, DUT.bus.q,
			);
		end
		T3: begin
			$display(
				"T3 @ %0t | PC=%0d MAR=%h MDR=%h IR=%h ALU_op=%0d Zlow=%0d reg_select=%b  R7=%h R0=%h R4=%h Y=%h Bus=%h",
				$time, DUT.PC.storage, DUT.MAR.storage, DUT.MDR.MDR_Reg.storage, DUT.IR.storage, ALU_operation, DUT.RZlow.storage, DUT.reg_decode, DUT.R7.storage, DUT.R0.storage, DUT.R4.storage, DUT.RY.storage, DUT.bus.q,
			);
		end
		T4: begin
			$display(
				"T4 @ %0t | PC=%0d MAR=%h MDR=%h IR=%h ALU_op=%0d Zlow=%0d reg_select=%b  R7=%h R0=%h R4=%h Y=%h Bus=%h",
				$time, DUT.PC.storage, DUT.MAR.storage, DUT.MDR.MDR_Reg.storage, DUT.IR.storage, ALU_operation, DUT.RZlow.storage, DUT.reg_decode, DUT.R7.storage, DUT.R0.storage, DUT.R4.storage, DUT.RY.storage, DUT.bus.q,
			);
		end
		T5: begin
			$display(
				"T5 @ %0t | PC=%0d MAR=%h MDR=%h IR=%h ALU_op=%0d Zlow=%0d reg_select=%b  R7=%h R0=%h R4=%h Y=%h Bus=%h",
				$time, DUT.PC.storage, DUT.MAR.storage, DUT.MDR.MDR_Reg.storage, DUT.IR.storage, ALU_operation, DUT.RZlow.storage, DUT.reg_decode, DUT.R7.storage, DUT.R0.storage, DUT.R4.storage, DUT.RY.storage, DUT.bus.q,
			);
		end
		done: begin
			$display(
				"End @ %0t | PC=%0d MAR=%h MDR=%h IR=%h ALU_op=%0d Zlow=%0d reg_select=%b R7=%h R0=%h R4=%h Y=%h Bus=%h",
				$time, DUT.PC.storage, DUT.MAR.storage, DUT.MDR.MDR_Reg.storage, DUT.IR.storage, ALU_operation, DUT.RZlow.storage, DUT.reg_decode, DUT.R7.storage, DUT.R0.storage, DUT.R4.storage, DUT.RY.storage, DUT.bus.q,
			);
			$stop;
		end
	endcase
end

endmodule 